module example2;
    int x, y, z;
    initial begin
        x = 1; y = 2; z = 3;
        $display("x: %d");
    end
endmodule
